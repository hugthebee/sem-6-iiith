
.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.global gnd vdd

Vdd	vdd	gnd	'SUPPLY'
vin a 0 pulse 0 1.8 0ns 1ns 1ns 10ns 20ns

.subckt inv y x vdd gnd
.param width_P={48*LAMBDA}
.param width_N={20*LAMBDA}
M1      y       x       gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
M2      y       x       vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
.ends inv

x1 b a vdd gnd inv
x2 c b vdd gnd inv

*.dc vin 0 1.8 0.1
.tran 0.1n 200n

** MEASURING DELAYS (Refer manual section 15.4.5)
.measure tran tperiod
+ TRIG v(b) VAL='SUPPLY/2' RISE=1
+ TARG v(b) VAL='SUPPLY/2' RISE=2
.measure tran tpdr
+ TRIG v(b) VAL='SUPPLY/2' FALL=1
+ TARG v(c) VAL='SUPPLY/2' RISE=1

.measure tran tpdf
+ TRIG v(b) VAL='SUPPLY/2' RISE=1
+ TARG v(c) VAL='SUPPLY/2' FALL=1

.measure tran tpd param='(tpdr+tpdf)/2' goal=0
.measure tran diff param='tpdr-tpdf' goal=0

.control
set hcopypscolor = 1 *White background for saving plots
set color0=white ** color0 is used to set the background of the plot (manual sec:17.7))
set color1=black ** color1 is used to set the grid color of the plot (manual sec:17.7))
set xbrushwidth = 3


run
*plot v(a)
*plot v(b)
plot  v(b) v(c)
plot i(vdd)

hardcopy fig_inv_trans.eps v(b) v(c)
.endc
